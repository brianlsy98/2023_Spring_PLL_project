** Generated for: hspiceD
** Generated on: May  6 15:14:42 2021
** Design library name: test
** Design cell name: osc
** Design view name: schematic


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: test
** Cell name: inv
** View name: schematic
.subckt inv in out vdd vss
m0 out in vss vss nmos L=45e-9 W=1e-6
m1 out in vdd vdd pmos L=45e-9 W=2e-6
.ends inv
** End of subcircuit definition.

** Library name: test
** Cell name: osc
** View name: schematic
xi11 net018 net031 vdd vss inv
xi10 net027 net029 vdd vss inv
xi8 net029 out vdd vss inv
xi7 net030 net027 vdd vss inv
xi6 net031 net030 vdd vss inv
xi5 net032 net034 vdd vss inv
xi4 net033 net018 vdd vss inv
xi3 net034 net033 vdd vss inv
xi2 net8 net032 vdd vss inv
xi1 net9 net8 vdd vss inv
xi0 out net9 vdd vss inv
.END
